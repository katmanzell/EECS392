
// I2C MPU-6050 Controller Module
// Usage: controls the 2-bus I2C module

// Clock is supposed to be at max i2c supported frequency!
	module top (
		clk,
		scl,
		sda,
		rst_n
);
	input clk;
	input	rst_n;
	output scl;
	output [7: 0] data;
	inout sda;

	reg [2: 0] cnt; // cnt = 0, rising scl; cnt = 1, scl high intermediate; cnt = 2, scl falling; cnt = 3, scl low intermediate
	reg [8: 0] cnt_sum; // generate the desired clock IIC
	reg scl_r; // clock pulse generated

	reg [19: 0] cnt_10ms;

	always @ (posedge clk or negedge rst_n)
	if (! rst_n)
	cnt_10ms <= 20'd0;
	else
	cnt_10ms <= cnt_10ms + 1'b1;

	always @ (posedge clk or negedge rst_n)
	begin
	if (! rst_n)
	cnt_sum <= 0;
	else if (cnt_sum == 9'd499)
	cnt_sum <= 0;
	else
	cnt_sum <= cnt_sum + 1'b1;
	end

	always @ (posedge clk or negedge rst_n)
	begin
	if (! rst_n)
	cnt <= 3'd5;
	else
	begin
	case (cnt_sum)
	9'd124: cnt <= 3'd1; // HIGH
	9'd249: cnt <= 3'd2; // falling
	9'd374: cnt <= 3'd3; // low
	9'd499: cnt <= 3'd0; // rising
	default: cnt <= 3'd5;
	endcase
	end
	end

	`Define SCL_POS (cnt == 3'd0);
	`Define SCL_HIG (cnt == 3'd1);
	`Define SCL_NEG (cnt == 3'd2);
	`Define SCL_LOW (cnt == 3'd3);

	always @ (posedge clk or negedge rst_n)
	begin
	if (! rst_n)
	scl_r <= 1'b0;
	else if (cnt == 3'd0)
	scl_r <= 1'b1;
	else if (cnt == 3'd2)
	scl_r <= 1'b0;
	end

	assign scl = scl_r; // scl clock signal

	`Define DEVICE_READ 8'hD1 // addressable device, read
	`Define DEVICE_WRITE 8'hD0 // addressable devices, writes
	`Define ACC_XH 8'h3B // x-axis acceleration upper address
	`Define ACC_XL 8'h3C // x-axis acceleration low address
	`Define ACC_YH 8'h3D // y-axis acceleration upper address
	`Define ACC_YL 8'h3E // y-axis acceleration low address
	`Define ACC_ZH 8'h3F // z axis acceleration upper address
	`Define ACC_ZL 8'h40 // z axis acceleration low address
	`Define GYRO_XH 8'h43 // x-axis gyroscope upper address
	`Define GYRO_XL 8'h44 // x-axis gyroscope low address
	`Define GYRO_YH 8'h45 // y-axis gyroscope upper address
	`Define GYRO_YL 8'h46 // y-axis gyroscope low address
	`Define GYRO_ZH 8'h47 // z-axis gyroscope upper address
	`Define GYRO_ZL 8'h48 // z-axis gyroscope low address

	// Initialize the registers gyroscope
	`Define PWR_MGMT_1 8'h6B
	`Define SMPLRT_DIV 8'h19
	`Define CONFIG1 8'h1A
	`Define GYRO_CONFIG 8'h1B
	`Define ACC_CONFIG 8'h1C
	// Gyroscope initialization value corresponds to the configuration register
	`Define PWR_MGMT_1_VAL 8'h00
	`Define SMPLRT_DIV_VAL 8'h07
	`Define CONFIG1_VAL 8'h06
	`Define GYRO_CONFIG_VAL 8'h18
	`Define ACC_CONFIG_VAL 8'h01

	parameter IDLE = 4'd0;
	parameter START1 = 4'd1;
	parameter ADD1 = 4'd2;
	parameter ACK1 = 4'd3;
	parameter ADD2 = 4'd4;
	parameter ACK2 = 4'd5;
	parameter START2 = 4'd6;
	parameter ADD3 = 4'd7;
	parameter ACK3 = 4'd8;
	parameter DATA = 4'd9;
	parameter ACK4 = 4'd10;
	parameter STOP1 = 4'd11;
	parameter STOP2 = 4'd12;
	parameter ADD_EXT = 4'd13;
	parameter ACK_EXT = 4'd14;

	reg [3: 0] state; // status register
	reg sda_r; // output
	reg sda_link; // sda_link = 1, sda output; sda_link = 0, sda high impedance
	reg [3: 0] num;
	reg [7: 0] db_r;
	reg [7: 0] ACC_XH_READ; // stored acceleration X-axis high eight
	reg [7: 0] ACC_XL_READ; // stored acceleration X-axis low eight
	reg [7: 0] ACC_YH_READ; // stored acceleration Y-axis high eight
	reg [7: 0] ACC_YL_READ; // low storage acceleration in the Y-axis eight
	reg [7: 0] ACC_ZH_READ; // stored acceleration Z axis high eight
	reg [7: 0] ACC_ZL_READ; // store the Z-axis acceleration low eight
	reg [7: 0] GYRO_XH_READ; // high storage X-axis gyroscope eight
	reg [7: 0] GYRO_XL_READ; // store low X-axis gyroscope eight
	reg [7: 0] GYRO_YH_READ; // store high Y-axis gyroscope eight
	reg [7: 0] GYRO_YL_READ; // Low memory Y-axis gyroscope eight
	reg [7: 0] GYRO_ZH_READ; // store gyroscope Z-axis high eight
	reg [7: 0] GYRO_ZL_READ; // store gyroscope Z-axis low eight
	reg [4: 0] times; // number of records initial configuration register

	always @ (posedge clk or negedge rst_n)
	begin
	if (! rst_n)
	begin
	state <= IDLE;
	sda_r <= 1'b1; // pulled data lines
	sda_link <= 1'b0; // high-impedance state
	num <= 4'd0;
	// Initialize the register
	ACC_XH_READ <= 8'h00;
	ACC_XL_READ <= 8'h00;
	ACC_YH_READ <= 8'h00;
	ACC_YL_READ <= 8'h00;
	ACC_ZH_READ <= 8'h00;
	ACC_ZL_READ <= 8'h00;
	GYRO_XH_READ <= 8'h00;
	GYRO_XL_READ <= 8'h00;
	GYRO_YH_READ <= 8'h00;
	GYRO_YL_READ <= 8'h00;
	GYRO_ZH_READ <= 8'h00;
	GYRO_ZL_READ <= 8'h00;
	times <= 5'b0;
	end
	else
	case (state)
	IDLE: begin
	times <= times + 1'b1;
	sda_link <= 1'b1; // sda output
	sda_r <= 1'b1; // pulled sda
	db_r <= `DEVICE_WRITE; // write data to the slave address
	state = START1;
	end
	START1: begin // IIC start
	if ( `SCL_HIG) // scl is high
	begin
	sda_link <= 1'b1; // sda output
	sda_r <= 1'b0; // low sda, generating start signal
	state <= ADD1;
	num <= 4'd0;
	end
	else
	state <= START1;
	end
	ADD1: begin // write data
	if ( `SCL_LOW) // scl low
	begin
	if (num == 4'd8) // When eight full output
	begin
	num <= 4'd0; // count is cleared
	sda_r <= 1'b1;
	sda_link <= 1'b0; // sda high impedance state
	state <= ACK1;
	end
	else
	begin
	state <= ADD1;
	num <= num + 1'b1;
	sda_r <= db_r [4'd7-num]; // bit output
	end
	end
	else
	state <= ADD1;
	end
	ACK1: begin // Answer
	if ( `SCL_NEG)
	begin
	state <= ADD2;
	case (times) // select the next write address register
	5'd1: db_r <= `PWR_MGMT_1;
	5'd2: db_r <= `SMPLRT_DIV;
	5'd3: db_r <= `CONFIG1;
	5'd4: db_r <= `GYRO_CONFIG;
	5'd5: db_r <= `ACC_CONFIG;
	5'd6: db_r <= `ACC_XH;
	5'd7: db_r <= `ACC_XL;
	5'd8: db_r <= `ACC_YH;
	5'd9: db_r <= `ACC_YL;
	5'd10: db_r <= `ACC_ZH;
	5'd11: db_r <= `ACC_ZL;
	5'd12: db_r <= `GYRO_XH;
	5'd13: db_r <= `GYRO_XL;
	5'd14: db_r <= `GYRO_YH;
	5'd15: db_r <= `GYRO_YL;
	5'd16: db_r <= `GYRO_ZH;
	5'd17: db_r <= `GYRO_ZL;
	default: begin
	db_r <= `PWR_MGMT_1;
	times <= 5'd1;
	end
	endcase
	end
	else
	state <= ACK1; // waits for a response
	end
	ADD2: begin
	if ( `SCL_LOW) // scl low
	begin
	if (num == 4'd8)
	begin
	num <= 4'd0;
	sda_r <= 1'b1;
	sda_link <= 1'b0;
	state <= ACK2;
	end
	else
	begin
	sda_link <= 1'b1;
	state <= ADD2;
	num <= num + 1'b1;
	sda_r <= db_r [4'd7-num]; // send bit address register
	end
	end
	else
	state <= ADD2;
	end
	ACK2: begin // Answer
	if ( `SCL_NEG)
	begin
	case (times) // set value of the corresponding register
	3'd1: db_r <= `PWR_MGMT_1_VAL;
	3'd2: db_r <= `SMPLRT_DIV_VAL;
	3'd3: db_r <= `CONFIG1_VAL;
	3'd4: db_r <= `GYRO_CONFIG_VAL;
	3'd5: db_r <= `ACC_CONFIG_VAL;
	3'd6: db_r <= `DEVICE_READ;
	default: db_r <= `DEVICE_READ;
	endcase
	if (times> = 5'd6)
	state <= START2;
	else
	state <= ADD_EXT;
	end
	else
	state <= ACK2; // waits for a response
	end
	ADD_EXT: begin // initialize some setting register
	if ( `SCL_LOW)
	begin
	if (num == 4'd8)
	begin
	num <= 4'd0;
	sda_r <= 1'b1;
	sda_link <= 1'b0; // sda high impedance state
	state <= ACK_EXT;
	end
	else
	begin
	sda_link <= 1'b1;
	state <= ADD_EXT;
	num <= num + 1'b1;
	sda_r <= db_r [4'd7-num]; // bit setting register work
	end
	end
	else
	state <= ADD_EXT;
	end
	ACK_EXT: begin
	if ( `SCL_NEG)
	begin
	sda_r <= 1'b1; // pulled sda
	state <= STOP1;
	end
	else
	state <= ACK_EXT; // waits for a response
	end
	START2: begin
	if ( `SCL_LOW) // scl low
	begin
	sda_link <= 1'b1; // sda output
	sda_r <= 1'b1; // pulled sda
	state <= START2;
	end
	else if ( `SCL_HIG) // scl is high
	begin
	sda_r <= 1'b0; // low sda, generating start signal
	state <= ADD3;
	end
	else
	state <= START2;
	end
	ADD3: begin
	if ( `SCL_LOW) // scl-bit low
	begin
	if (num == 4'd8)
	begin
	num <= 4'd0;
	sda_r <= 1'b1; // pulled sda
	sda_link <= 1'b0; // scl high impedance state
	state <= ACK3;
	end
	else
	begin
	num <= num + 1'b1;
	sda_r <= db_r [4'd7-num]; // write bit read register address
	state <= ADD3;
	end
	end
	else state <= ADD3;
	end
	ACK3: begin
	if ( `SCL_NEG)
	begin
	state <= DATA;
	sda_link <= 1'b0; // sda high impedance state
	end
	else
	state <= ACK3; // waits for a response
	end
	DATA: begin
	if (num <= 4'd7)
	begin
	state <= DATA;
	if ( `SCL_HIG)
	begin
	num <= num + 1'b1;
	case (times)
	5'd6: ACC_XH_READ [4'd7-num] <= sda;
	5'd7: ACC_XL_READ [4'd7-num] <= sda;
	5'd8: ACC_YH_READ [4'd7-num] <= sda;
	5'd9: ACC_YL_READ [4'd7-num] <= sda;
	5'd10: ACC_ZH_READ [4'd7-num] <= sda;
	5'd11: ACC_ZL_READ [4'd7-num] <= sda;
	5'd12: GYRO_XH_READ [4'd7-num] <= sda;
	5'd13: GYRO_XL_READ [4'd7-num] <= sda;
	5'd14: GYRO_YH_READ [4'd7-num] <= sda;
	5'd15: GYRO_YL_READ [4'd7-num] <= sda;
	5'd16: GYRO_ZH_READ [4'd7-num] <= sda;
	5'd17: GYRO_ZL_READ [4'd7-num] <= sda;
	default:; // not yet considered, can add code to improve system stability
	endcase
	end
	end
	else if (( `SCL_LOW) && (num == 4'd8))
	begin
	sda_link <= 1'b1; // sda output
	num <= 4'd0; // count is cleared
	state <= ACK4;
	end
	else
	state <= DATA;
	end
	ACK4: begin
	if (times == 5'd17)
	times <= 5'd0;
	if ( `SCL_NEG)
	begin
	sda_r <= 1'b1; // pulled sda
	state <= STOP1;
	end
	else
	state <= ACK4; // waits for a response
	end
	STOP1: begin
	if ( `SCL_LOW) // scl low
	begin
	sda_link <= 1'b1; // sda output
	sda_r <= 1'b0; // low sda
	state <= STOP1;
	end
	else if ( `SCL_HIG) // sda high
	begin
	sda_r <= 1'b1; // pulled sda, generates stop signal
	state <= STOP2;
	end
	else
	state <= STOP1;
	end
	STOP2: begin
	if ( `SCL_LOW)
	sda_r <= 1'b1;
	else if (cnt_10ms == 20'hffff0) // get data about 10ms
	state <= IDLE;
	else
	state <= STOP2;
	end
	default: state <= IDLE;
	endcase
	end

	assign sda = sda_link sda_r: 1'bz;?

	endmodule